module instr_mem
(  
	input			[15:0]	pc,  
	output wire	[15:0]	instruction  
);  

	wire [3:0] rom_addr = pc[3:0];

	/* 
	lw $3, 0($0) --   
	Loop: slti $1, $3, 50  
	beq $1, $0, Skip  
	add $4, $4, $3   
	addi $3, $3, 1   
	beq $0, $0, Loop--  
	Skip  
	*/

	reg [15:0] rom[15:0];  
	
	initial  
	begin  
	
		rom[0]	= 16'h444f;
		rom[1]	= 16'h465f;
		rom[2]	= 16'h14c0;
		rom[3]	= 16'h0000;
		rom[4]	= 16'h0000;
		rom[5]	= 16'h0000;
		rom[6]	= 16'h0000;
		rom[7]	= 16'h0000;  
		rom[8]	= 16'h0000;  
		rom[9]	= 16'h0000;  
		rom[10]	= 16'h0000;  
		rom[11]	= 16'h0000;
		rom[12]	= 16'h0000;  
		rom[13]	= 16'h0000;  
		rom[14]	= 16'h0000;  
		rom[15]	= 16'h0000;  
	
	end  
	
	assign instruction = (pc[15:0] < 16) ? rom[ rom_addr[3:0] ] : 16'd0;

endmodule